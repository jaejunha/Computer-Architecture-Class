
module Datapath(clk, reset_n);
	input clk;
	input reset_n;
endmodule